** Library name: work_VR
** Cell name: tgate
** View name: schematic

.subckt tgate in out vdda vssa

m0 in  vdda out vssa nch L=180e-9 W=1.8e-6 M=1
m1 out vssa in  vdda pch L=180e-9 W=4.0e-6 M=2

.ends tgate
** End of subcircuit definition.
