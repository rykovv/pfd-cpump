** Library name: work_VR
** Cell name: inverter
** View name: schematic

.subckt inverter in out vdda vssa

m0 out in vdda vdda pch L=180e-9 W=4.0e-6 M=2
m1 out in vssa vssa nch L=180e-9 W=1.8e-6 M=1

.ends inverter
** End of subcircuit definition.
